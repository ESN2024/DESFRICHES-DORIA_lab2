
module counter (
	clk_clk,
	reset_reset_n,
	pio_0_external_connection_export);	

	input		clk_clk;
	input		reset_reset_n;
	output	[3:0]	pio_0_external_connection_export;
endmodule
